// === defines.sv ===
 
`define IV_0 32'h6A09E667
`define IV_1 32'hBB67AE85
`define IV_2 32'h3C6EF372
`define IV_3 32'hA54FF53A
`define IV_4 32'h510e527f
`define IV_5 32'h9b05688c
`define IV_6 32'h1f83d9ab
`define IV_7 32'h5be0cd19
